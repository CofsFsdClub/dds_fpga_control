`define SUPPORT_RV32C 1
`define SUPPORT_RV32M 1
`define ENABLE_COUNTERS 1
`define ENABLE_IRQ 1
`define ENABLE_TIMER 1
`define TWO_STAGE_SHIFT 1
`define TWO_CYCLE_COMPARE 0
`define TWO_CYCLE_ALU 0
`define BARREL_SHIFTER 0
`define CATCH_MISALIGN 1
`define CATCH_ILLINSN 1
`define ENABLE_DEBUG
`define I_MEM_K_BYTE 64
`define BUILD_LOAD
`define SW_BIN_PATH "D:/Program_Station/Embedded_Program/GOWIN_FPGA/dds_project/mcu_projecct/Debug/ram32.hex"
`define D_MEM_K_BYTE 32
`define ENABLE_HSP 0
`define HSP_VALUE_DEF 32'h0
`define ENABLE_WB_GPIO
`define GPIO_DW 4
`define ENABLE_ADVSPI
`define ADVSPI_REG
`define ADVSPI_MEM_SUPPORT
`define ENABLE_SIMPLE_UART
`define ENABLE_WB_UART
`define ENABLE_WB_SPI_MASTER
`define WBSPI_MASTER_SHIFT_DIRECTION 0
`define WBSPI_MASTER_CLOCK_PHASE 0
`define WBSPI_MASTER_CLOCK_POLARITY 0
`define WBSPI_MASTER_CLKCNT_WIDTH 10
`define WBSPI_MASTER_CLOCK_SEL 2
`define WBSPI_MASTER_SLAVE_NUMBER 1
`define WBSPI_MASTER_DATA_LENGTH 8
`define WBSPI_MASTER_DELAY_TIME 1
`define WBSPI_MASTER_INTERVAL_LENGTH 1
`define DEVICE_ARORA_V
